* G:\Users\richa_000\Google Drive 2\Sous Vide Files\Hardware\SousVide.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 28/09/2017 16:49:25

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ATMEGA328PB-AU		
U2  ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? Net-_U2-Pad33_ Net-_U2-Pad33_ Net-_U2-Pad33_ Net-_U2-Pad36_ Net-_U2-Pad36_ Net-_U2-Pad36_ MAX6954		
U3  ? ? /O0 ? ? ? ? /O0 ? ? 7SEGMENT_CC		
U5  ? ? /O1 ? ? ? ? /O1 ? ? 7SEGMENT_CC		
U4  ? ? /O2 ? ? ? ? /O2 ? ? 7SEGMENT_CC		
U6  ? ? /O3 ? ? ? ? /O3 ? ? 7SEGMENT_CC		

.end
